`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   01:45:19 02/28/2015
// Design Name:   cache_test
// Module Name:   C:/Users/lgonza20/Desktop/lab4/lab4/sim_cache_test.v
// Project Name:  lab4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: cache_test
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module sim_cache_test;

	// Inputs
	reg clk;
	reg rst;
	reg we;
	reg [31:0] mem_data;
	reg rd;
	reg [31:0] addr;

	// Outputs
	wire [31:0] mem_addr;
	wire valid;
	wire [31:0] data;
	//wire [31:0] reg_addr;
	wire hit,miss;
	wire [2:0] way;
	wire [23:0] tag,tag_check;
	wire [1:0] lru1,lru2,lru3,lru4;
	wire [5:0] state;

	// Instantiate the Unit Under Test (UUT)
	cache_test uut (
		.clk(clk), 
		.rst(rst), 
		.we(we), 
		.mem_data(mem_data), 
		.mem_addr(mem_addr), 
		.rd(rd), 
		.addr(addr), 
		.valid(valid), 
		.data(data),
		//.reg_addr(reg_addr),
		.hit(hit),
		.miss(miss),
		.way(way),
		.tag(tag),
		.tag_check(tag_check),
		.lru1(lru1),
		.lru2(lru2),
		.lru3(lru3),
		.lru4(lru4),
		
		.state(state)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		we = 0;
		mem_data = 0;
		rd = 0;
		addr = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'hFFFF_DC00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		mem_data <= 32'h ABCD_0000;
		#5
		clk=1;
		we=1;
		mem_data <= 32'h ABCD_0000;
		#5
		clk=0;
		#5
		clk=1;
		mem_data <= 32'h0000_0000;
		we=0;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'hDDDD_DD00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr =32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'hCCCC_CC00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		mem_data = 32'h5678_5678;
		#5
		clk=1;
		we=1;
		mem_data = 32'h5678_5678;
		#5
		clk=0;
		#5
		clk=1;
		we=0;
		mem_data = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'hFFFF_FF00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'h8888_8800;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		mem_data=32'h1234_1234;
		#5
		clk=1;
		we=1;
		mem_data=32'h1234_1234;
		#5
		clk=0;
		#5
		clk=1;
		we=0;
		mem_data=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		//addr = 32'hDDDD_DD00;
		addr=32'hCCCC_CC00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		//addr=32'hCCCC_CC00;
		addr = 32'hDDDD_DD00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		mem_data=32'h1111_1111;
		#5
		clk=1;
		we=1;
		mem_data=32'h1111_1111;
		#5
		clk=0;
		#5
		clk=1;
		we=0;
		mem_data=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'habcd_0000;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'h1111_1100;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		

	end
      
endmodule

