`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:12:23 02/24/2015 
// Design Name: 
// Module Name:    compare 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//module compare(input clk,
//					input [31:0] addr_reg,
//					input [23:0] tag,
//					output result
//    );
//	 
//	 always @(*)begin
//		if(tag==addr_reg[31:7]) // assuming tag is 24 bits
//			results = 1'b1;
//		else
//			result = 1'b0;
//	end
//	
//	 
//	 
//
//
//endmodule
