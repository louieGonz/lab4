`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:30:25 02/24/2015
// Design Name:   block
// Module Name:   C:/Users/lgonza20/Desktop/lab4/lab4/sim_block.v
// Project Name:  lab4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: block
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module sim_block;

	// Inputs
	reg clk;
	reg rd;
	reg [31:0] addr;
	
	

	// Outputs
	wire hit;
	wire [31:0] reg_addr;
	wire [23:0] tag;
	wire [23:0] tag_check;
	wire [2:0] way;
	wire miss;
	wire atMM;
	wire [4:0] state;
	wire [1:0] outMM;
	wire [1:0] way1set0;
	wire [1:0] way2set0;
	wire [1:0] way3set0;
	wire [1:0] way4set0;
	wire [31:0] way1data,way2data,way3data,way4data;

	// Instantiate the Unit Under Test (UUT)
	block uut (
		.clk(clk),
		.rd(rd),
		.addr(addr),
		.reg_addr(reg_addr),
		.tag(tag),
		.tag_check(tag_check),
		.way(way),
		.miss(miss),
		.atMM(atMM),
		.state(state),
		.outMM(outMM),
		.way1set0(way1set0),
		.way2set0(way2set0),
		.way3set0(way3set0),
		.way4set0(way4set0),
		.way1data(way1data),
		.way2data(way2data),
		.way3data(way3data),
		.way4data(way4data),
		.hit(hit)
	);

	initial begin
		// Initialize Inputs
		clk = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		//addr =  32'h0000_0000;
		#5
		clk=1;
		//rd=1;
		//addr = 32'hFFFF_FF00;
		#5
		clk=0;
		#5
		clk=1;
		//addr = 32'h0000_0000;
		rd=0;
		
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr =  32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		#5
		clk=0;
		#5
		clk=1;
		//rd=0;
		#5
		clk=0;
		#5
		clk=1;
		//rd=1;
		//addr = 32'hFFFF_FF;
		#5
		clk=0;
		#5
		clk=1;
		//addr = 32'h0000_0000;
		//rd=0;
		#5
		clk=0;
		#5
		clk=1;
		//rd=1;
		//addr =  32'h0000_0003;
		#5
		clk=0;
		#5
		clk=1;
		//rd=0;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		//addr = 32'hFFFF_FFF5;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'hFFFF_FF00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'h0000_ABC2;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'hCCCC_CC00;
		#5
		clk=0;
		#5
		rd=0;
		addr =32'h0000_0000;
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'h3333_3300;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'hDDDD_DD00;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr=32'h0000_0100;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr=32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		rd=1;
		addr = 32'h0000_00FD;
		#5
		clk=0;
		#5
		clk=1;
		rd=0;
		addr = 32'h0000_0000;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		#5
		clk=1;
		#5
		clk=0;
		


	end
      
endmodule

